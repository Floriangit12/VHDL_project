Création capteur moteur
